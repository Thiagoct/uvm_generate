interface xxx_if
	(
		input logic clk,
		input logic rst
	);

endinterface 	